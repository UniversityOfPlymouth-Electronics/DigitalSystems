module parity_challenge #(parameter N=8) (output logic P, input logic [N-1:0] X);


endmodule



