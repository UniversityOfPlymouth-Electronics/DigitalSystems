module mux2_structural (output logic y, input logic a, b, s);

// Write HDL here


endmodule