module pressrelease_tb_solution;

